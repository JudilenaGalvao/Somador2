library verilog;
use verilog.vl_types.all;
entity somador2_vlg_vec_tst is
end somador2_vlg_vec_tst;
